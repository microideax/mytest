`define FEATURE_WIDTH 8    //(include 1bit sign)

`define KERNEL_SIZE 5
`define KERNEL_WIDTH 2     //ternary complement -1 0 1 



`define IMAGE_IN_BIT_WIDTH 8
`define IMAGE_IN_WIDTH 32
`define IMAGE_IN_HEIGHT 32

